* AD8017 Spice Macro-model
* Description: Amplifier
* Generic Desc: Dual high speed 16dBm output op amp
* Developed by: JCH/CentApps
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (01/1999)
* Copyright 1999, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*
* Parameters modeled include:
*
* END Notes
*
* Node assignments
*                non-inverting input
*                |  inverting input
*                |  |  positive supply
*                |  |  |  negative supply
*                |  |  |  |  output
*                |  |  |  |  |
.SUBCKT AD8017   +I -1 +V -V Vo


***** Input Stage

q1   4  4 41 qn1
q2   3  3 41 qp1
i1  99  4 1.5e-4
i2   3 50 1.5e-4
cin1 1 88 2.4pf
q3   9 4 2 qn2
q4  10 3 2 qp2

rxxa  99  4 100k
rxxb   3 50 100k

VT1    9 99 0
VT2   10 50 0

vos   41  1 1.8m
fnoi1  1  0 vn2 1
fnoi2  2  0 vn2 1

***** internal inoise source

vbi 73 88 0.545
dn2 73 72 dninv
rn3 72 88 36
vn2 72 88 0

***** internal reference

Eref 88 0 poly(2) 99 0 50 0 0 0.5 0.5

***** gain stage/dominant pole/clamp circuitry

F3  29 88 VT1 1
F4  29 88 VT2 1
r3  29 88 710k
c1  29 88 1.84p

vc1 99 45 1.59
vc2 46 50 1.59
dc1 29 45 dx
dc2 46 29 dx

***** pole at 177MHz

egain2 32 88 88 29 1
r4     32 44 1
c3     44 88 0.835n

***** buffer to output stage

gbuf 34 88 44 88 1e-2
re1  34 88 100

***** output stage

fo1   88 110 vcd 1
do1  110 111 dx
do2  112 110 dx
vi1  111  88 0
vi2   88 112 0

fsy1  99  0 poly(2) visy1 vi1 6.3e-3 -1 1
fsy2   0 50 poly(2) visy2 vi2 6.3e-3 -1 1

go3   60 63 99 34 2.5
go4   64 60 34 50 2.5
r03   60 63 0.4
r04   60 64 0.4
visy1 99 63 0
visy2 64 50 0
vcd   60 61 0
do5   34 70 dx
do6   71 34 dx
vo1   70 60 -0.405
vo2   60 71 -0.405

.model dx d(is=1e-13 kf=6.5e-20 af=0)
.model dninv d(kf=5e-14)
.model qn1 npn(bf=200)
.model qn2 npn(bf=200)
.model qp1 pnp(bf=200)
.model qp2 pnp(bf=200)
.ends ad8017





